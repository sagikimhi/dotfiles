//-----------------------------------------------------------------------------
// Project       : Pixie
//-----------------------------------------------------------------------------
//
// File          : env_module.svh
// Author        : sagikimhi
// Created       : Thu Mar 2025, 23:10:47
// Last modified : Thu Mar 2025, 23:10:47
//
//-----------------------------------------------------------------------------
// Copyright (c) Wiliot.
//------------------------------------------------------------------------------
// Modification history:
// Thu Mar 2025, 23:10:47
//-----------------------------------------------------------------------------

`ifndef ENV_MODULE_SVH
`define ENV_MODULE_SVH

`timescale 1ns / 1ps

`include "uvm_macros.h"

module env_module
    import uvm_pkg::*;
#(
    parameter uvm_active_passive_enum ACTIVE_PASSIVE = uvm_pkg::UVM_ACTIVE
)
(
    input logic clk,
    input logic rst_n
);

    // ---------------------------------------------------------------------------
    // Wire Declarations
    // ---------------------------------------------------------------------------

    // ---------------------------------------------------------------------------
    // Interface Declarations
    // ---------------------------------------------------------------------------

    // ---------------------------------------------------------------------------
    // Interface Conntections
    // ---------------------------------------------------------------------------

    generate
    endgenerate

    // ---------------------------------------------------------------------------
    // Run Test
    // ---------------------------------------------------------------------------

    initial begin
        uvm_pkg::run_test();
        $finish();
    end

endmodule: env_module

`endif // ENV_MODULE_SVH
